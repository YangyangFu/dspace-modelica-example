<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<Root>
	<creator type="key">ConfigurationDesk 6.5</creator>
	<application>
		<Name type="key">ModelicaConstant.CDL</Name>
		<DisplayName type="key">ModelicaConstant</DisplayName>
		<Path type="key">.\ModelicaConstant</Path>
		<Component type="key">ProjectApplication</Component>
		<Type type="key">14</Type>
		<ApplicationType type="key">3</ApplicationType>
		<Flags type="key">41216</Flags>
		<ItemInfoDate type="key">10/6/2021 2:28:43 PM</ItemInfoDate>
		<ItemInfoPath type="key">$FPATH$</ItemInfoPath>
		<ItemInfoDocs type="key"/>
		<ItemInfoDescr type="key"/>
		<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
		<Log type="key"/>
		<AddInfoDb type="key"/>
		<DatabaseID type="key">-1</DatabaseID>
		<EntityID type="key">{B6725FDA-87B8-4C13-9826-C9F863A29945}</EntityID>
		<item>
			<Name type="key">WindowConfiguration.xml</Name>
			<DisplayName type="key">WindowConfiguration.xml</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">260</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">4</Type>
			<ItemInfoDate type="key">10/8/2021 4:56:20 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{8A6B08FA-C0DF-4A00-81E1-5221675580A0}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Device Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">33</Type>
			<ItemInfoDate type="key">10/6/2021 2:28:46 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{DEBB76B7-A049-4DC4-8DDB-CB792F5106CB}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Hardware Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">19</Type>
			<ItemInfoDate type="key">10/6/2021 2:28:46 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{6F7FA835-FECF-4D06-BAB0-AAB5B29C7B70}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Model Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">31</Type>
			<ItemInfoDate type="key">10/6/2021 2:28:46 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key">Model location:
D:\github\dspace-modelica-example\dSpaceExample\ds_modelica_constant.slx
</Log>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{5B1625BF-54A1-4396-A4C6-178A942BB732}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Communication Matrices</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">70</Type>
			<ItemInfoDate type="key">10/6/2021 2:28:46 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{96B93E3D-E1D3-4A27-AD83-E851445CEEA5}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">External Cable Harness</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">32</Type>
			<ItemInfoDate type="key">10/6/2021 2:28:46 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{564B4953-C012-4421-B6F4-4CAA4C557278}</EntityID>
			<Targets/>
		</item>
		<item>
			<Name type="key">Application.cfgx</Name>
			<DisplayName type="key">Core Application</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">260</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">20</Type>
			<ItemInfoDate type="key">10/6/2021 2:28:46 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{BC48FAF3-6521-4434-9E73-15E0C3EBDFBD}</EntityID>
			<Targets/>
		</item>
		<item>
			<Name type="key">Build Results</Name>
			<DisplayName type="key">Build Results</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">58</Type>
			<ItemInfoDate type="key">10/8/2021 4:57:37 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{41935818-7D0A-46B5-9D01-145FD0E87D3C}</EntityID>
			<Targets/>
			<item>
				<Name type="key">Build Results</Name>
				<DisplayName type="key">itSDFROOT</DisplayName>
				<Path type="key">.</Path>
				<Component type="key">ProjectApplication</Component>
				<Flags type="key">260</Flags>
				<ExtendedFlags type="key">0</ExtendedFlags>
				<Type type="key">29</Type>
				<ItemInfoDate type="key">10/8/2021 4:57:37 PM</ItemInfoDate>
				<ItemInfoPath type="key"/>
				<ItemInfoDocs type="key"/>
				<ItemInfoDescr type="key"/>
				<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
				<ItemInfoAddInfoDb type="key"/>
				<Log type="key"/>
				<DatabaseID type="key">-1</DatabaseID>
				<EntityID type="key">{B382A75B-102D-4C66-93AC-EADDAB7D0CAA}</EntityID>
				<Targets/>
				<item>
					<Name type="key">ds_modelica_constant.expswcfg</Name>
					<DisplayName type="key">ds_modelica_constant.expswcfg</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">71</Type>
					<ItemInfoDate type="key">10/8/2021 4:57:37 PM</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{572B691C-C321-49BC-B579-A4B4E630803D}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">ds_modelica_constant.map</Name>
					<DisplayName type="key">ds_modelica_constant.map</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">36</Type>
					<ItemInfoDate type="key">10/8/2021 4:57:37 PM</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{BC1C4D5B-EAE5-4588-A70A-9DE528B50CED}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">ds_modelica_constant.trc</Name>
					<DisplayName type="key">ds_modelica_constant.trc</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">34</Type>
					<ItemInfoDate type="key">10/8/2021 4:57:37 PM</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{C9DF5A37-F039-4C3F-97DD-FD04E53750B3}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">ModelicaConstant.dsbuildinfo</Name>
					<DisplayName type="key">ModelicaConstant.dsbuildinfo</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">260</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">4</Type>
					<ItemInfoDate type="key">10/8/2021 4:57:37 PM</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{9D6CECF4-5100-41AD-A51B-F3D0770DD862}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">ModelicaConstant.rta</Name>
					<DisplayName type="key">ModelicaConstant.rta</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">37</Type>
					<ItemInfoDate type="key">10/8/2021 4:57:37 PM</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{9701B5C7-BF05-4F94-A769-FDF7E3BF625F}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">ModelicaConstant.sdf</Name>
					<DisplayName type="key">ModelicaConstant.sdf</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">35</Type>
					<ItemInfoDate type="key">10/8/2021 4:57:37 PM</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{D8AFF52A-12E2-4B73-8C74-32FE0458D4FC}</EntityID>
					<Targets/>
				</item>
			</item>
		</item>
	</application>
</Root>