<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<Root>
	<creator type="key">ConfigurationDesk 6.5</creator>
	<application>
		<Name type="key">twozone_outputs.CDL</Name>
		<DisplayName type="key">twozone_outputs</DisplayName>
		<Path type="key">.\twozone_outputs</Path>
		<Component type="key">ProjectApplication</Component>
		<Type type="key">14</Type>
		<ApplicationType type="key">3</ApplicationType>
		<Flags type="key">41216</Flags>
		<ItemInfoDate type="key">9/29/2021 6:06:13 PM</ItemInfoDate>
		<ItemInfoPath type="key">$FPATH$</ItemInfoPath>
		<ItemInfoDocs type="key"/>
		<ItemInfoDescr type="key"/>
		<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
		<Log type="key"/>
		<AddInfoDb type="key"/>
		<DatabaseID type="key">-1</DatabaseID>
		<EntityID type="key">{A5B48817-FBB7-42F8-9378-1C101E9709E7}</EntityID>
		<item>
			<Name type="key">WindowConfiguration.xml</Name>
			<DisplayName type="key">WindowConfiguration.xml</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">260</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">4</Type>
			<ItemInfoDate type="key">10/6/2021 2:15:04 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{1F079914-7512-4EAB-8C05-6F6F3FB22769}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Device Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">33</Type>
			<ItemInfoDate type="key">9/29/2021 6:06:15 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{903EE1B6-0EF9-4F58-88AB-B4AAE48D3282}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Hardware Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">19</Type>
			<ItemInfoDate type="key">9/29/2021 6:06:15 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{CCE80EB2-6432-48D9-943C-1BC4B98F45E2}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Model Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">31</Type>
			<ItemInfoDate type="key">9/29/2021 6:06:15 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key">Model location:
D:\github\dspace-modelica-example\dSpaceExample\ds_fivezoneg36_dsrt.slx
</Log>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{49B78E1A-1195-4668-AA70-DF4CE66F8BFA}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Communication Matrices</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">70</Type>
			<ItemInfoDate type="key">9/29/2021 6:06:15 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{8E49EE3D-7933-4D64-9805-BA371C9D3650}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">External Cable Harness</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">32</Type>
			<ItemInfoDate type="key">9/29/2021 6:06:15 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{D303B586-1669-494C-A2C2-AAE82146AC07}</EntityID>
			<Targets/>
		</item>
		<item>
			<Name type="key">Application.cfgx</Name>
			<DisplayName type="key">Core Application</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">260</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">20</Type>
			<ItemInfoDate type="key">9/29/2021 6:06:15 PM</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">yangyang.fu</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{CE811EAD-4811-43A3-8DBD-32D2274744BB}</EntityID>
			<Targets/>
		</item>
	</application>
</Root>